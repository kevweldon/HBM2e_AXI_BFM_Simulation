// my_sys.v

// Generated using ACDS version 22.4 94

`timescale 1 ps / 1 ps
module my_sys (
		input  wire       axi_reset_in_reset,                      //          axi_reset_in.reset
		input  wire       clk100_in_clk,                           //             clk100_in.clk
		input  wire       hbm_reset_in_reset,                      //          hbm_reset_in.reset
		input  wire       hbm_fp_0_cattrip_i_conduit,              //    hbm_fp_0_cattrip_i.conduit
		input  wire [2:0] hbm_fp_0_temp_i_conduit,                 //       hbm_fp_0_temp_i.conduit
		output wire       hbm_local_cal_success_local_cal_success, // hbm_local_cal_success.local_cal_success
		output wire       hbm_local_cal_fail_local_cal_fail,       //    hbm_local_cal_fail.local_cal_fail
		output wire       hbm_wmcrst_n_reset_n,                    //          hbm_wmcrst_n.reset_n
		output wire       iopll_locked_export,                     //          iopll_locked.export
		input  wire       iopll_reset_reset,                       //           iopll_reset.reset
		input  wire       noc_reset_in_reset                       //          noc_reset_in.reset
	);

	wire          clk100_out_clk_clk;                                      // clk100:out_clk -> [intel_noc_clock_ctrl_0:refclk, iopll_0:refclk]
	wire          iopll_0_outclk0_clk;                                     // iopll_0:outclk_0 -> [intel_noc_initiator_0:s_axi4_aclk, mgc_axi4_master_0:ACLK, mgc_axi4_master_1:ACLK, mm_interconnect_0:iopll_0_outclk0_clk, mm_interconnect_1:iopll_0_outclk0_clk, rst_controller:clk, rst_controller_001:clk, rst_controller_002:clk]
	wire          iopll_0_outclk1_clk;                                     // iopll_0:outclk_1 -> hbm_fp_0:uibpll_refclk
	wire          noc_reset_out_reset_reset;                               // noc_reset:out_reset -> [intel_noc_initiator_0:s_axi4_aresetn, rst_controller_002:reset_in0]
	wire    [7:0] mgc_axi4_master_0_altera_axi4_master_ruser;              // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_ruser -> mgc_axi4_master_0:RUSER
	wire    [7:0] mgc_axi4_master_0_altera_axi4_master_wuser;              // mgc_axi4_master_0:WUSER -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_wuser
	wire    [1:0] mgc_axi4_master_0_altera_axi4_master_awburst;            // mgc_axi4_master_0:AWBURST -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awburst
	wire    [3:0] mgc_axi4_master_0_altera_axi4_master_arregion;           // mgc_axi4_master_0:ARREGION -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arregion
	wire    [7:0] mgc_axi4_master_0_altera_axi4_master_arlen;              // mgc_axi4_master_0:ARLEN -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arlen
	wire    [3:0] mgc_axi4_master_0_altera_axi4_master_arqos;              // mgc_axi4_master_0:ARQOS -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arqos
	wire    [7:0] mgc_axi4_master_0_altera_axi4_master_awuser;             // mgc_axi4_master_0:AWUSER -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awuser
	wire          mgc_axi4_master_0_altera_axi4_master_wready;             // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_wready -> mgc_axi4_master_0:WREADY
	wire   [31:0] mgc_axi4_master_0_altera_axi4_master_wstrb;              // mgc_axi4_master_0:WSTRB -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_wstrb
	wire    [6:0] mgc_axi4_master_0_altera_axi4_master_rid;                // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_rid -> mgc_axi4_master_0:RID
	wire          mgc_axi4_master_0_altera_axi4_master_rready;             // mgc_axi4_master_0:RREADY -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_rready
	wire    [7:0] mgc_axi4_master_0_altera_axi4_master_awlen;              // mgc_axi4_master_0:AWLEN -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awlen
	wire    [3:0] mgc_axi4_master_0_altera_axi4_master_awqos;              // mgc_axi4_master_0:AWQOS -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awqos
	wire          mgc_axi4_master_0_altera_axi4_master_wvalid;             // mgc_axi4_master_0:WVALID -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_wvalid
	wire   [63:0] mgc_axi4_master_0_altera_axi4_master_araddr;             // mgc_axi4_master_0:ARADDR -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_araddr
	wire    [2:0] mgc_axi4_master_0_altera_axi4_master_arprot;             // mgc_axi4_master_0:ARPROT -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arprot
	wire    [2:0] mgc_axi4_master_0_altera_axi4_master_awprot;             // mgc_axi4_master_0:AWPROT -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awprot
	wire          mgc_axi4_master_0_altera_axi4_master_arvalid;            // mgc_axi4_master_0:ARVALID -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arvalid
	wire  [255:0] mgc_axi4_master_0_altera_axi4_master_wdata;              // mgc_axi4_master_0:WDATA -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_wdata
	wire    [6:0] mgc_axi4_master_0_altera_axi4_master_arid;               // mgc_axi4_master_0:ARID -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arid
	wire          mgc_axi4_master_0_altera_axi4_master_arlock;             // mgc_axi4_master_0:ARLOCK -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arlock
	wire          mgc_axi4_master_0_altera_axi4_master_awlock;             // mgc_axi4_master_0:AWLOCK -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awlock
	wire   [63:0] mgc_axi4_master_0_altera_axi4_master_awaddr;             // mgc_axi4_master_0:AWADDR -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awaddr
	wire          mgc_axi4_master_0_altera_axi4_master_arready;            // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arready -> mgc_axi4_master_0:ARREADY
	wire    [1:0] mgc_axi4_master_0_altera_axi4_master_bresp;              // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_bresp -> mgc_axi4_master_0:BRESP
	wire  [255:0] mgc_axi4_master_0_altera_axi4_master_rdata;              // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_rdata -> mgc_axi4_master_0:RDATA
	wire          mgc_axi4_master_0_altera_axi4_master_awready;            // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awready -> mgc_axi4_master_0:AWREADY
	wire    [1:0] mgc_axi4_master_0_altera_axi4_master_arburst;            // mgc_axi4_master_0:ARBURST -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arburst
	wire    [2:0] mgc_axi4_master_0_altera_axi4_master_arsize;             // mgc_axi4_master_0:ARSIZE -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_arsize
	wire          mgc_axi4_master_0_altera_axi4_master_rlast;              // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_rlast -> mgc_axi4_master_0:RLAST
	wire          mgc_axi4_master_0_altera_axi4_master_bready;             // mgc_axi4_master_0:BREADY -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_bready
	wire          mgc_axi4_master_0_altera_axi4_master_wlast;              // mgc_axi4_master_0:WLAST -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_wlast
	wire    [3:0] mgc_axi4_master_0_altera_axi4_master_awregion;           // mgc_axi4_master_0:AWREGION -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awregion
	wire    [1:0] mgc_axi4_master_0_altera_axi4_master_rresp;              // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_rresp -> mgc_axi4_master_0:RRESP
	wire    [6:0] mgc_axi4_master_0_altera_axi4_master_awid;               // mgc_axi4_master_0:AWID -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awid
	wire    [6:0] mgc_axi4_master_0_altera_axi4_master_bid;                // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_bid -> mgc_axi4_master_0:BID
	wire          mgc_axi4_master_0_altera_axi4_master_bvalid;             // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_bvalid -> mgc_axi4_master_0:BVALID
	wire          mgc_axi4_master_0_altera_axi4_master_awvalid;            // mgc_axi4_master_0:AWVALID -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awvalid
	wire    [2:0] mgc_axi4_master_0_altera_axi4_master_awsize;             // mgc_axi4_master_0:AWSIZE -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_awsize
	wire          mgc_axi4_master_0_altera_axi4_master_rvalid;             // mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_rvalid -> mgc_axi4_master_0:RVALID
	wire    [7:0] mgc_axi4_master_0_altera_axi4_master_aruser;             // mgc_axi4_master_0:ARUSER -> mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_aruser
	wire   [31:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_ruser;   // intel_noc_initiator_0:s0_axi4_ruser -> mm_interconnect_0:intel_noc_initiator_0_s0_axi4_ruser
	wire   [31:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wuser;   // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_wuser -> intel_noc_initiator_0:s0_axi4_wuser
	wire    [1:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awburst; // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_awburst -> intel_noc_initiator_0:s0_axi4_awburst
	wire   [10:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awuser;  // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_awuser -> intel_noc_initiator_0:s0_axi4_awuser
	wire    [7:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arlen;   // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_arlen -> intel_noc_initiator_0:s0_axi4_arlen
	wire    [3:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arqos;   // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_arqos -> intel_noc_initiator_0:s0_axi4_arqos
	wire   [31:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wstrb;   // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_wstrb -> intel_noc_initiator_0:s0_axi4_wstrb
	wire          mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wready;  // intel_noc_initiator_0:s0_axi4_wready -> mm_interconnect_0:intel_noc_initiator_0_s0_axi4_wready
	wire    [6:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rid;     // intel_noc_initiator_0:s0_axi4_rid -> mm_interconnect_0:intel_noc_initiator_0_s0_axi4_rid
	wire          mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rready;  // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_rready -> intel_noc_initiator_0:s0_axi4_rready
	wire    [7:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awlen;   // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_awlen -> intel_noc_initiator_0:s0_axi4_awlen
	wire    [3:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awqos;   // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_awqos -> intel_noc_initiator_0:s0_axi4_awqos
	wire          mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wvalid;  // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_wvalid -> intel_noc_initiator_0:s0_axi4_wvalid
	wire   [43:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_araddr;  // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_araddr -> intel_noc_initiator_0:s0_axi4_araddr
	wire    [2:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arprot;  // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_arprot -> intel_noc_initiator_0:s0_axi4_arprot
	wire    [2:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awprot;  // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_awprot -> intel_noc_initiator_0:s0_axi4_awprot
	wire  [255:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wdata;   // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_wdata -> intel_noc_initiator_0:s0_axi4_wdata
	wire          mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arvalid; // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_arvalid -> intel_noc_initiator_0:s0_axi4_arvalid
	wire    [6:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arid;    // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_arid -> intel_noc_initiator_0:s0_axi4_arid
	wire    [0:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arlock;  // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_arlock -> intel_noc_initiator_0:s0_axi4_arlock
	wire    [0:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awlock;  // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_awlock -> intel_noc_initiator_0:s0_axi4_awlock
	wire   [43:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awaddr;  // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_awaddr -> intel_noc_initiator_0:s0_axi4_awaddr
	wire    [1:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_bresp;   // intel_noc_initiator_0:s0_axi4_bresp -> mm_interconnect_0:intel_noc_initiator_0_s0_axi4_bresp
	wire          mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arready; // intel_noc_initiator_0:s0_axi4_arready -> mm_interconnect_0:intel_noc_initiator_0_s0_axi4_arready
	wire  [255:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rdata;   // intel_noc_initiator_0:s0_axi4_rdata -> mm_interconnect_0:intel_noc_initiator_0_s0_axi4_rdata
	wire          mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awready; // intel_noc_initiator_0:s0_axi4_awready -> mm_interconnect_0:intel_noc_initiator_0_s0_axi4_awready
	wire    [1:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arburst; // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_arburst -> intel_noc_initiator_0:s0_axi4_arburst
	wire    [2:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arsize;  // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_arsize -> intel_noc_initiator_0:s0_axi4_arsize
	wire          mm_interconnect_0_intel_noc_initiator_0_s0_axi4_bready;  // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_bready -> intel_noc_initiator_0:s0_axi4_bready
	wire          mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rlast;   // intel_noc_initiator_0:s0_axi4_rlast -> mm_interconnect_0:intel_noc_initiator_0_s0_axi4_rlast
	wire          mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wlast;   // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_wlast -> intel_noc_initiator_0:s0_axi4_wlast
	wire    [1:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rresp;   // intel_noc_initiator_0:s0_axi4_rresp -> mm_interconnect_0:intel_noc_initiator_0_s0_axi4_rresp
	wire    [6:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awid;    // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_awid -> intel_noc_initiator_0:s0_axi4_awid
	wire    [6:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_bid;     // intel_noc_initiator_0:s0_axi4_bid -> mm_interconnect_0:intel_noc_initiator_0_s0_axi4_bid
	wire          mm_interconnect_0_intel_noc_initiator_0_s0_axi4_bvalid;  // intel_noc_initiator_0:s0_axi4_bvalid -> mm_interconnect_0:intel_noc_initiator_0_s0_axi4_bvalid
	wire    [2:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awsize;  // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_awsize -> intel_noc_initiator_0:s0_axi4_awsize
	wire          mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awvalid; // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_awvalid -> intel_noc_initiator_0:s0_axi4_awvalid
	wire   [10:0] mm_interconnect_0_intel_noc_initiator_0_s0_axi4_aruser;  // mm_interconnect_0:intel_noc_initiator_0_s0_axi4_aruser -> intel_noc_initiator_0:s0_axi4_aruser
	wire          mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rvalid;  // intel_noc_initiator_0:s0_axi4_rvalid -> mm_interconnect_0:intel_noc_initiator_0_s0_axi4_rvalid
	wire    [7:0] mgc_axi4_master_1_altera_axi4_master_ruser;              // mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_ruser -> mgc_axi4_master_1:RUSER
	wire    [7:0] mgc_axi4_master_1_altera_axi4_master_wuser;              // mgc_axi4_master_1:WUSER -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_wuser
	wire    [1:0] mgc_axi4_master_1_altera_axi4_master_awburst;            // mgc_axi4_master_1:AWBURST -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_awburst
	wire    [3:0] mgc_axi4_master_1_altera_axi4_master_arregion;           // mgc_axi4_master_1:ARREGION -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_arregion
	wire    [7:0] mgc_axi4_master_1_altera_axi4_master_arlen;              // mgc_axi4_master_1:ARLEN -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_arlen
	wire    [3:0] mgc_axi4_master_1_altera_axi4_master_arqos;              // mgc_axi4_master_1:ARQOS -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_arqos
	wire    [7:0] mgc_axi4_master_1_altera_axi4_master_awuser;             // mgc_axi4_master_1:AWUSER -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_awuser
	wire          mgc_axi4_master_1_altera_axi4_master_wready;             // mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_wready -> mgc_axi4_master_1:WREADY
	wire   [31:0] mgc_axi4_master_1_altera_axi4_master_wstrb;              // mgc_axi4_master_1:WSTRB -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_wstrb
	wire    [6:0] mgc_axi4_master_1_altera_axi4_master_rid;                // mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_rid -> mgc_axi4_master_1:RID
	wire          mgc_axi4_master_1_altera_axi4_master_rready;             // mgc_axi4_master_1:RREADY -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_rready
	wire    [7:0] mgc_axi4_master_1_altera_axi4_master_awlen;              // mgc_axi4_master_1:AWLEN -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_awlen
	wire    [3:0] mgc_axi4_master_1_altera_axi4_master_awqos;              // mgc_axi4_master_1:AWQOS -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_awqos
	wire          mgc_axi4_master_1_altera_axi4_master_wvalid;             // mgc_axi4_master_1:WVALID -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_wvalid
	wire   [63:0] mgc_axi4_master_1_altera_axi4_master_araddr;             // mgc_axi4_master_1:ARADDR -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_araddr
	wire    [2:0] mgc_axi4_master_1_altera_axi4_master_arprot;             // mgc_axi4_master_1:ARPROT -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_arprot
	wire    [2:0] mgc_axi4_master_1_altera_axi4_master_awprot;             // mgc_axi4_master_1:AWPROT -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_awprot
	wire          mgc_axi4_master_1_altera_axi4_master_arvalid;            // mgc_axi4_master_1:ARVALID -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_arvalid
	wire  [255:0] mgc_axi4_master_1_altera_axi4_master_wdata;              // mgc_axi4_master_1:WDATA -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_wdata
	wire    [6:0] mgc_axi4_master_1_altera_axi4_master_arid;               // mgc_axi4_master_1:ARID -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_arid
	wire          mgc_axi4_master_1_altera_axi4_master_arlock;             // mgc_axi4_master_1:ARLOCK -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_arlock
	wire          mgc_axi4_master_1_altera_axi4_master_awlock;             // mgc_axi4_master_1:AWLOCK -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_awlock
	wire   [63:0] mgc_axi4_master_1_altera_axi4_master_awaddr;             // mgc_axi4_master_1:AWADDR -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_awaddr
	wire          mgc_axi4_master_1_altera_axi4_master_arready;            // mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_arready -> mgc_axi4_master_1:ARREADY
	wire    [1:0] mgc_axi4_master_1_altera_axi4_master_bresp;              // mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_bresp -> mgc_axi4_master_1:BRESP
	wire  [255:0] mgc_axi4_master_1_altera_axi4_master_rdata;              // mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_rdata -> mgc_axi4_master_1:RDATA
	wire          mgc_axi4_master_1_altera_axi4_master_awready;            // mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_awready -> mgc_axi4_master_1:AWREADY
	wire    [1:0] mgc_axi4_master_1_altera_axi4_master_arburst;            // mgc_axi4_master_1:ARBURST -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_arburst
	wire    [2:0] mgc_axi4_master_1_altera_axi4_master_arsize;             // mgc_axi4_master_1:ARSIZE -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_arsize
	wire          mgc_axi4_master_1_altera_axi4_master_rlast;              // mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_rlast -> mgc_axi4_master_1:RLAST
	wire          mgc_axi4_master_1_altera_axi4_master_bready;             // mgc_axi4_master_1:BREADY -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_bready
	wire          mgc_axi4_master_1_altera_axi4_master_wlast;              // mgc_axi4_master_1:WLAST -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_wlast
	wire    [3:0] mgc_axi4_master_1_altera_axi4_master_awregion;           // mgc_axi4_master_1:AWREGION -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_awregion
	wire    [1:0] mgc_axi4_master_1_altera_axi4_master_rresp;              // mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_rresp -> mgc_axi4_master_1:RRESP
	wire    [6:0] mgc_axi4_master_1_altera_axi4_master_awid;               // mgc_axi4_master_1:AWID -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_awid
	wire    [6:0] mgc_axi4_master_1_altera_axi4_master_bid;                // mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_bid -> mgc_axi4_master_1:BID
	wire          mgc_axi4_master_1_altera_axi4_master_bvalid;             // mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_bvalid -> mgc_axi4_master_1:BVALID
	wire          mgc_axi4_master_1_altera_axi4_master_awvalid;            // mgc_axi4_master_1:AWVALID -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_awvalid
	wire    [2:0] mgc_axi4_master_1_altera_axi4_master_awsize;             // mgc_axi4_master_1:AWSIZE -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_awsize
	wire          mgc_axi4_master_1_altera_axi4_master_rvalid;             // mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_rvalid -> mgc_axi4_master_1:RVALID
	wire    [7:0] mgc_axi4_master_1_altera_axi4_master_aruser;             // mgc_axi4_master_1:ARUSER -> mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_aruser
	wire   [31:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_ruser;   // intel_noc_initiator_0:s1_axi4_ruser -> mm_interconnect_1:intel_noc_initiator_0_s1_axi4_ruser
	wire   [31:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wuser;   // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_wuser -> intel_noc_initiator_0:s1_axi4_wuser
	wire    [1:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awburst; // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_awburst -> intel_noc_initiator_0:s1_axi4_awburst
	wire   [10:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awuser;  // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_awuser -> intel_noc_initiator_0:s1_axi4_awuser
	wire    [7:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arlen;   // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_arlen -> intel_noc_initiator_0:s1_axi4_arlen
	wire    [3:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arqos;   // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_arqos -> intel_noc_initiator_0:s1_axi4_arqos
	wire   [31:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wstrb;   // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_wstrb -> intel_noc_initiator_0:s1_axi4_wstrb
	wire          mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wready;  // intel_noc_initiator_0:s1_axi4_wready -> mm_interconnect_1:intel_noc_initiator_0_s1_axi4_wready
	wire    [6:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rid;     // intel_noc_initiator_0:s1_axi4_rid -> mm_interconnect_1:intel_noc_initiator_0_s1_axi4_rid
	wire          mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rready;  // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_rready -> intel_noc_initiator_0:s1_axi4_rready
	wire    [7:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awlen;   // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_awlen -> intel_noc_initiator_0:s1_axi4_awlen
	wire    [3:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awqos;   // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_awqos -> intel_noc_initiator_0:s1_axi4_awqos
	wire          mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wvalid;  // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_wvalid -> intel_noc_initiator_0:s1_axi4_wvalid
	wire   [43:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_araddr;  // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_araddr -> intel_noc_initiator_0:s1_axi4_araddr
	wire    [2:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arprot;  // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_arprot -> intel_noc_initiator_0:s1_axi4_arprot
	wire    [2:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awprot;  // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_awprot -> intel_noc_initiator_0:s1_axi4_awprot
	wire  [255:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wdata;   // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_wdata -> intel_noc_initiator_0:s1_axi4_wdata
	wire          mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arvalid; // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_arvalid -> intel_noc_initiator_0:s1_axi4_arvalid
	wire    [6:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arid;    // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_arid -> intel_noc_initiator_0:s1_axi4_arid
	wire    [0:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arlock;  // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_arlock -> intel_noc_initiator_0:s1_axi4_arlock
	wire    [0:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awlock;  // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_awlock -> intel_noc_initiator_0:s1_axi4_awlock
	wire   [43:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awaddr;  // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_awaddr -> intel_noc_initiator_0:s1_axi4_awaddr
	wire    [1:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_bresp;   // intel_noc_initiator_0:s1_axi4_bresp -> mm_interconnect_1:intel_noc_initiator_0_s1_axi4_bresp
	wire          mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arready; // intel_noc_initiator_0:s1_axi4_arready -> mm_interconnect_1:intel_noc_initiator_0_s1_axi4_arready
	wire  [255:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rdata;   // intel_noc_initiator_0:s1_axi4_rdata -> mm_interconnect_1:intel_noc_initiator_0_s1_axi4_rdata
	wire          mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awready; // intel_noc_initiator_0:s1_axi4_awready -> mm_interconnect_1:intel_noc_initiator_0_s1_axi4_awready
	wire    [1:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arburst; // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_arburst -> intel_noc_initiator_0:s1_axi4_arburst
	wire    [2:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arsize;  // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_arsize -> intel_noc_initiator_0:s1_axi4_arsize
	wire          mm_interconnect_1_intel_noc_initiator_0_s1_axi4_bready;  // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_bready -> intel_noc_initiator_0:s1_axi4_bready
	wire          mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rlast;   // intel_noc_initiator_0:s1_axi4_rlast -> mm_interconnect_1:intel_noc_initiator_0_s1_axi4_rlast
	wire          mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wlast;   // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_wlast -> intel_noc_initiator_0:s1_axi4_wlast
	wire    [1:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rresp;   // intel_noc_initiator_0:s1_axi4_rresp -> mm_interconnect_1:intel_noc_initiator_0_s1_axi4_rresp
	wire    [6:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awid;    // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_awid -> intel_noc_initiator_0:s1_axi4_awid
	wire    [6:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_bid;     // intel_noc_initiator_0:s1_axi4_bid -> mm_interconnect_1:intel_noc_initiator_0_s1_axi4_bid
	wire          mm_interconnect_1_intel_noc_initiator_0_s1_axi4_bvalid;  // intel_noc_initiator_0:s1_axi4_bvalid -> mm_interconnect_1:intel_noc_initiator_0_s1_axi4_bvalid
	wire    [2:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awsize;  // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_awsize -> intel_noc_initiator_0:s1_axi4_awsize
	wire          mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awvalid; // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_awvalid -> intel_noc_initiator_0:s1_axi4_awvalid
	wire   [10:0] mm_interconnect_1_intel_noc_initiator_0_s1_axi4_aruser;  // mm_interconnect_1:intel_noc_initiator_0_s1_axi4_aruser -> intel_noc_initiator_0:s1_axi4_aruser
	wire          mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rvalid;  // intel_noc_initiator_0:s1_axi4_rvalid -> mm_interconnect_1:intel_noc_initiator_0_s1_axi4_rvalid
	wire          rst_controller_reset_out_reset;                          // rst_controller:reset_out -> [mgc_axi4_master_0:ARESETn, mgc_axi4_master_1:ARESETn]
	wire          axi_reset_out_reset_reset;                               // axi_reset:out_reset -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	wire          rst_controller_001_reset_out_reset;                      // rst_controller_001:reset_out -> [mm_interconnect_0:mgc_axi4_master_0_altera_axi4_master_translator_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:mgc_axi4_master_1_altera_axi4_master_translator_clk_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_002_reset_out_reset;                      // rst_controller_002:reset_out -> [mm_interconnect_0:intel_noc_initiator_0_s0_axi4_translator_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_1:intel_noc_initiator_0_s1_axi4_translator_clk_reset_reset_bridge_in_reset_reset]

	axi_reset axi_reset (
		.in_reset  (axi_reset_in_reset),        //   input,  width = 1,  in_reset.reset
		.out_reset (axi_reset_out_reset_reset)  //  output,  width = 1, out_reset.reset
	);

	clk100 clk100 (
		.in_clk  (clk100_in_clk),      //   input,  width = 1,  in_clk.clk
		.out_clk (clk100_out_clk_clk)  //  output,  width = 1, out_clk.clk
	);

	my_sys_hbm_fp_0 hbm_fp_0 (
		.ch0_u0_wmc_intr   (),                                        //  output,  width = 1,   ch0_u0_wmc_intr.conduit
		.ch0_u1_wmc_intr   (),                                        //  output,  width = 1,   ch0_u1_wmc_intr.conduit
		.hbm_reset_in      (hbm_reset_in_reset),                      //   input,  width = 1,      hbm_reset_in.reset
		.hbm_cattrip       (),                                        //  output,  width = 1,           cattrip.hbm_cattrip
		.hbm_cattrip_i     (hbm_fp_0_cattrip_i_conduit),              //   input,  width = 1,         cattrip_i.conduit
		.hbm_temp          (),                                        //  output,  width = 3,              temp.hbm_temp
		.hbm_temp_i        (hbm_fp_0_temp_i_conduit),                 //   input,  width = 3,            temp_i.conduit
		.local_cal_success (hbm_local_cal_success_local_cal_success), //  output,  width = 1, local_cal_success.local_cal_success
		.local_cal_fail    (hbm_local_cal_fail_local_cal_fail),       //  output,  width = 1,    local_cal_fail.local_cal_fail
		.uibpll_refclk     (iopll_0_outclk1_clk),                     //   input,  width = 1,     uibpll_refclk.clk
		.wmcrst_n          (hbm_wmcrst_n_reset_n)                     //  output,  width = 1,          wmcrst_n.reset_n
	);

	my_sys_intel_noc_clock_ctrl_0 intel_noc_clock_ctrl_0 (
		.refclk     (clk100_out_clk_clk), //   input,  width = 1,     refclk.clk
		.pll_lock_o ()                    //  output,  width = 1, pll_lock_o.pll_lock_o
	);

	my_sys_intel_noc_initiator_0 intel_noc_initiator_0 (
		.s0_axi4_awid    (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awid),    //   input,    width = 7,        s0_axi4.awid
		.s0_axi4_awaddr  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awaddr),  //   input,   width = 44,               .awaddr
		.s0_axi4_awlen   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awlen),   //   input,    width = 8,               .awlen
		.s0_axi4_awsize  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awsize),  //   input,    width = 3,               .awsize
		.s0_axi4_awburst (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awburst), //   input,    width = 2,               .awburst
		.s0_axi4_awlock  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awlock),  //   input,    width = 1,               .awlock
		.s0_axi4_awprot  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awprot),  //   input,    width = 3,               .awprot
		.s0_axi4_awuser  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awuser),  //   input,   width = 11,               .awuser
		.s0_axi4_awqos   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awqos),   //   input,    width = 4,               .awqos
		.s0_axi4_awvalid (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awvalid), //   input,    width = 1,               .awvalid
		.s0_axi4_awready (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awready), //  output,    width = 1,               .awready
		.s0_axi4_wdata   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wdata),   //   input,  width = 256,               .wdata
		.s0_axi4_wstrb   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wstrb),   //   input,   width = 32,               .wstrb
		.s0_axi4_wlast   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wlast),   //   input,    width = 1,               .wlast
		.s0_axi4_wvalid  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wvalid),  //   input,    width = 1,               .wvalid
		.s0_axi4_wuser   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wuser),   //   input,   width = 32,               .wuser
		.s0_axi4_wready  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wready),  //  output,    width = 1,               .wready
		.s0_axi4_bid     (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_bid),     //  output,    width = 7,               .bid
		.s0_axi4_bresp   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_bresp),   //  output,    width = 2,               .bresp
		.s0_axi4_bvalid  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_bvalid),  //  output,    width = 1,               .bvalid
		.s0_axi4_bready  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_bready),  //   input,    width = 1,               .bready
		.s0_axi4_arid    (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arid),    //   input,    width = 7,               .arid
		.s0_axi4_araddr  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_araddr),  //   input,   width = 44,               .araddr
		.s0_axi4_arlen   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arlen),   //   input,    width = 8,               .arlen
		.s0_axi4_arsize  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arsize),  //   input,    width = 3,               .arsize
		.s0_axi4_arburst (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arburst), //   input,    width = 2,               .arburst
		.s0_axi4_arlock  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arlock),  //   input,    width = 1,               .arlock
		.s0_axi4_arprot  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arprot),  //   input,    width = 3,               .arprot
		.s0_axi4_aruser  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_aruser),  //   input,   width = 11,               .aruser
		.s0_axi4_arqos   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arqos),   //   input,    width = 4,               .arqos
		.s0_axi4_arvalid (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arvalid), //   input,    width = 1,               .arvalid
		.s0_axi4_arready (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arready), //  output,    width = 1,               .arready
		.s0_axi4_rid     (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rid),     //  output,    width = 7,               .rid
		.s0_axi4_rdata   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rdata),   //  output,  width = 256,               .rdata
		.s0_axi4_rresp   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rresp),   //  output,    width = 2,               .rresp
		.s0_axi4_rlast   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rlast),   //  output,    width = 1,               .rlast
		.s0_axi4_rvalid  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rvalid),  //  output,    width = 1,               .rvalid
		.s0_axi4_rready  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rready),  //   input,    width = 1,               .rready
		.s0_axi4_ruser   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_ruser),   //  output,   width = 32,               .ruser
		.s1_axi4_awid    (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awid),    //   input,    width = 7,        s1_axi4.awid
		.s1_axi4_awaddr  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awaddr),  //   input,   width = 44,               .awaddr
		.s1_axi4_awlen   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awlen),   //   input,    width = 8,               .awlen
		.s1_axi4_awsize  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awsize),  //   input,    width = 3,               .awsize
		.s1_axi4_awburst (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awburst), //   input,    width = 2,               .awburst
		.s1_axi4_awlock  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awlock),  //   input,    width = 1,               .awlock
		.s1_axi4_awprot  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awprot),  //   input,    width = 3,               .awprot
		.s1_axi4_awuser  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awuser),  //   input,   width = 11,               .awuser
		.s1_axi4_awqos   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awqos),   //   input,    width = 4,               .awqos
		.s1_axi4_awvalid (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awvalid), //   input,    width = 1,               .awvalid
		.s1_axi4_awready (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awready), //  output,    width = 1,               .awready
		.s1_axi4_wdata   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wdata),   //   input,  width = 256,               .wdata
		.s1_axi4_wstrb   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wstrb),   //   input,   width = 32,               .wstrb
		.s1_axi4_wlast   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wlast),   //   input,    width = 1,               .wlast
		.s1_axi4_wvalid  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wvalid),  //   input,    width = 1,               .wvalid
		.s1_axi4_wuser   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wuser),   //   input,   width = 32,               .wuser
		.s1_axi4_wready  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wready),  //  output,    width = 1,               .wready
		.s1_axi4_bid     (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_bid),     //  output,    width = 7,               .bid
		.s1_axi4_bresp   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_bresp),   //  output,    width = 2,               .bresp
		.s1_axi4_bvalid  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_bvalid),  //  output,    width = 1,               .bvalid
		.s1_axi4_bready  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_bready),  //   input,    width = 1,               .bready
		.s1_axi4_arid    (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arid),    //   input,    width = 7,               .arid
		.s1_axi4_araddr  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_araddr),  //   input,   width = 44,               .araddr
		.s1_axi4_arlen   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arlen),   //   input,    width = 8,               .arlen
		.s1_axi4_arsize  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arsize),  //   input,    width = 3,               .arsize
		.s1_axi4_arburst (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arburst), //   input,    width = 2,               .arburst
		.s1_axi4_arlock  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arlock),  //   input,    width = 1,               .arlock
		.s1_axi4_arprot  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arprot),  //   input,    width = 3,               .arprot
		.s1_axi4_aruser  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_aruser),  //   input,   width = 11,               .aruser
		.s1_axi4_arqos   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arqos),   //   input,    width = 4,               .arqos
		.s1_axi4_arvalid (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arvalid), //   input,    width = 1,               .arvalid
		.s1_axi4_arready (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arready), //  output,    width = 1,               .arready
		.s1_axi4_rid     (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rid),     //  output,    width = 7,               .rid
		.s1_axi4_rdata   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rdata),   //  output,  width = 256,               .rdata
		.s1_axi4_rresp   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rresp),   //  output,    width = 2,               .rresp
		.s1_axi4_rlast   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rlast),   //  output,    width = 1,               .rlast
		.s1_axi4_rvalid  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rvalid),  //  output,    width = 1,               .rvalid
		.s1_axi4_rready  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rready),  //   input,    width = 1,               .rready
		.s1_axi4_ruser   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_ruser),   //  output,   width = 32,               .ruser
		.s_axi4_aclk     (iopll_0_outclk0_clk),                                     //   input,    width = 1,    s_axi4_aclk.clk
		.s_axi4_aresetn  (~noc_reset_out_reset_reset)                               //   input,    width = 1, s_axi4_aresetn.reset_n
	);

	my_sys_iopll_0 iopll_0 (
		.refclk   (clk100_out_clk_clk),  //   input,  width = 1,  refclk.clk
		.locked   (iopll_locked_export), //  output,  width = 1,  locked.export
		.rst      (iopll_reset_reset),   //   input,  width = 1,   reset.reset
		.outclk_0 (iopll_0_outclk0_clk), //  output,  width = 1, outclk0.clk
		.outclk_1 (iopll_0_outclk1_clk)  //  output,  width = 1, outclk1.clk
	);

	my_sys_mgc_axi4_master_0 mgc_axi4_master_0 (
		.AWVALID  (mgc_axi4_master_0_altera_axi4_master_awvalid),  //  output,    width = 1, altera_axi4_master.awvalid
		.AWPROT   (mgc_axi4_master_0_altera_axi4_master_awprot),   //  output,    width = 3,                   .awprot
		.AWREGION (mgc_axi4_master_0_altera_axi4_master_awregion), //  output,    width = 4,                   .awregion
		.AWLEN    (mgc_axi4_master_0_altera_axi4_master_awlen),    //  output,    width = 8,                   .awlen
		.AWSIZE   (mgc_axi4_master_0_altera_axi4_master_awsize),   //  output,    width = 3,                   .awsize
		.AWBURST  (mgc_axi4_master_0_altera_axi4_master_awburst),  //  output,    width = 2,                   .awburst
		.AWLOCK   (mgc_axi4_master_0_altera_axi4_master_awlock),   //  output,    width = 1,                   .awlock
		.AWQOS    (mgc_axi4_master_0_altera_axi4_master_awqos),    //  output,    width = 4,                   .awqos
		.AWREADY  (mgc_axi4_master_0_altera_axi4_master_awready),  //   input,    width = 1,                   .awready
		.ARVALID  (mgc_axi4_master_0_altera_axi4_master_arvalid),  //  output,    width = 1,                   .arvalid
		.ARPROT   (mgc_axi4_master_0_altera_axi4_master_arprot),   //  output,    width = 3,                   .arprot
		.ARREGION (mgc_axi4_master_0_altera_axi4_master_arregion), //  output,    width = 4,                   .arregion
		.ARLEN    (mgc_axi4_master_0_altera_axi4_master_arlen),    //  output,    width = 8,                   .arlen
		.ARSIZE   (mgc_axi4_master_0_altera_axi4_master_arsize),   //  output,    width = 3,                   .arsize
		.ARBURST  (mgc_axi4_master_0_altera_axi4_master_arburst),  //  output,    width = 2,                   .arburst
		.ARLOCK   (mgc_axi4_master_0_altera_axi4_master_arlock),   //  output,    width = 1,                   .arlock
		.ARQOS    (mgc_axi4_master_0_altera_axi4_master_arqos),    //  output,    width = 4,                   .arqos
		.ARREADY  (mgc_axi4_master_0_altera_axi4_master_arready),  //   input,    width = 1,                   .arready
		.RVALID   (mgc_axi4_master_0_altera_axi4_master_rvalid),   //   input,    width = 1,                   .rvalid
		.RRESP    (mgc_axi4_master_0_altera_axi4_master_rresp),    //   input,    width = 2,                   .rresp
		.RLAST    (mgc_axi4_master_0_altera_axi4_master_rlast),    //   input,    width = 1,                   .rlast
		.RREADY   (mgc_axi4_master_0_altera_axi4_master_rready),   //  output,    width = 1,                   .rready
		.WVALID   (mgc_axi4_master_0_altera_axi4_master_wvalid),   //  output,    width = 1,                   .wvalid
		.WLAST    (mgc_axi4_master_0_altera_axi4_master_wlast),    //  output,    width = 1,                   .wlast
		.WREADY   (mgc_axi4_master_0_altera_axi4_master_wready),   //   input,    width = 1,                   .wready
		.BVALID   (mgc_axi4_master_0_altera_axi4_master_bvalid),   //   input,    width = 1,                   .bvalid
		.BRESP    (mgc_axi4_master_0_altera_axi4_master_bresp),    //   input,    width = 2,                   .bresp
		.BREADY   (mgc_axi4_master_0_altera_axi4_master_bready),   //  output,    width = 1,                   .bready
		.AWADDR   (mgc_axi4_master_0_altera_axi4_master_awaddr),   //  output,   width = 64,                   .awaddr
		.AWID     (mgc_axi4_master_0_altera_axi4_master_awid),     //  output,    width = 7,                   .awid
		.AWUSER   (mgc_axi4_master_0_altera_axi4_master_awuser),   //  output,    width = 8,                   .awuser
		.ARADDR   (mgc_axi4_master_0_altera_axi4_master_araddr),   //  output,   width = 64,                   .araddr
		.ARID     (mgc_axi4_master_0_altera_axi4_master_arid),     //  output,    width = 7,                   .arid
		.ARUSER   (mgc_axi4_master_0_altera_axi4_master_aruser),   //  output,    width = 8,                   .aruser
		.RUSER    (mgc_axi4_master_0_altera_axi4_master_ruser),    //   input,    width = 8,                   .ruser
		.WUSER    (mgc_axi4_master_0_altera_axi4_master_wuser),    //  output,    width = 8,                   .wuser
		.RDATA    (mgc_axi4_master_0_altera_axi4_master_rdata),    //   input,  width = 256,                   .rdata
		.RID      (mgc_axi4_master_0_altera_axi4_master_rid),      //   input,    width = 7,                   .rid
		.WDATA    (mgc_axi4_master_0_altera_axi4_master_wdata),    //  output,  width = 256,                   .wdata
		.WSTRB    (mgc_axi4_master_0_altera_axi4_master_wstrb),    //  output,   width = 32,                   .wstrb
		.BID      (mgc_axi4_master_0_altera_axi4_master_bid),      //   input,    width = 7,                   .bid
		.ACLK     (iopll_0_outclk0_clk),                           //   input,    width = 1,         clock_sink.clk
		.ARESETn  (~rst_controller_reset_out_reset)                //   input,    width = 1,         reset_sink.reset_n
	);

	my_sys_mgc_axi4_master_0 mgc_axi4_master_1 (
		.AWVALID  (mgc_axi4_master_1_altera_axi4_master_awvalid),  //  output,    width = 1, altera_axi4_master.awvalid
		.AWPROT   (mgc_axi4_master_1_altera_axi4_master_awprot),   //  output,    width = 3,                   .awprot
		.AWREGION (mgc_axi4_master_1_altera_axi4_master_awregion), //  output,    width = 4,                   .awregion
		.AWLEN    (mgc_axi4_master_1_altera_axi4_master_awlen),    //  output,    width = 8,                   .awlen
		.AWSIZE   (mgc_axi4_master_1_altera_axi4_master_awsize),   //  output,    width = 3,                   .awsize
		.AWBURST  (mgc_axi4_master_1_altera_axi4_master_awburst),  //  output,    width = 2,                   .awburst
		.AWLOCK   (mgc_axi4_master_1_altera_axi4_master_awlock),   //  output,    width = 1,                   .awlock
		.AWQOS    (mgc_axi4_master_1_altera_axi4_master_awqos),    //  output,    width = 4,                   .awqos
		.AWREADY  (mgc_axi4_master_1_altera_axi4_master_awready),  //   input,    width = 1,                   .awready
		.ARVALID  (mgc_axi4_master_1_altera_axi4_master_arvalid),  //  output,    width = 1,                   .arvalid
		.ARPROT   (mgc_axi4_master_1_altera_axi4_master_arprot),   //  output,    width = 3,                   .arprot
		.ARREGION (mgc_axi4_master_1_altera_axi4_master_arregion), //  output,    width = 4,                   .arregion
		.ARLEN    (mgc_axi4_master_1_altera_axi4_master_arlen),    //  output,    width = 8,                   .arlen
		.ARSIZE   (mgc_axi4_master_1_altera_axi4_master_arsize),   //  output,    width = 3,                   .arsize
		.ARBURST  (mgc_axi4_master_1_altera_axi4_master_arburst),  //  output,    width = 2,                   .arburst
		.ARLOCK   (mgc_axi4_master_1_altera_axi4_master_arlock),   //  output,    width = 1,                   .arlock
		.ARQOS    (mgc_axi4_master_1_altera_axi4_master_arqos),    //  output,    width = 4,                   .arqos
		.ARREADY  (mgc_axi4_master_1_altera_axi4_master_arready),  //   input,    width = 1,                   .arready
		.RVALID   (mgc_axi4_master_1_altera_axi4_master_rvalid),   //   input,    width = 1,                   .rvalid
		.RRESP    (mgc_axi4_master_1_altera_axi4_master_rresp),    //   input,    width = 2,                   .rresp
		.RLAST    (mgc_axi4_master_1_altera_axi4_master_rlast),    //   input,    width = 1,                   .rlast
		.RREADY   (mgc_axi4_master_1_altera_axi4_master_rready),   //  output,    width = 1,                   .rready
		.WVALID   (mgc_axi4_master_1_altera_axi4_master_wvalid),   //  output,    width = 1,                   .wvalid
		.WLAST    (mgc_axi4_master_1_altera_axi4_master_wlast),    //  output,    width = 1,                   .wlast
		.WREADY   (mgc_axi4_master_1_altera_axi4_master_wready),   //   input,    width = 1,                   .wready
		.BVALID   (mgc_axi4_master_1_altera_axi4_master_bvalid),   //   input,    width = 1,                   .bvalid
		.BRESP    (mgc_axi4_master_1_altera_axi4_master_bresp),    //   input,    width = 2,                   .bresp
		.BREADY   (mgc_axi4_master_1_altera_axi4_master_bready),   //  output,    width = 1,                   .bready
		.AWADDR   (mgc_axi4_master_1_altera_axi4_master_awaddr),   //  output,   width = 64,                   .awaddr
		.AWID     (mgc_axi4_master_1_altera_axi4_master_awid),     //  output,    width = 7,                   .awid
		.AWUSER   (mgc_axi4_master_1_altera_axi4_master_awuser),   //  output,    width = 8,                   .awuser
		.ARADDR   (mgc_axi4_master_1_altera_axi4_master_araddr),   //  output,   width = 64,                   .araddr
		.ARID     (mgc_axi4_master_1_altera_axi4_master_arid),     //  output,    width = 7,                   .arid
		.ARUSER   (mgc_axi4_master_1_altera_axi4_master_aruser),   //  output,    width = 8,                   .aruser
		.RUSER    (mgc_axi4_master_1_altera_axi4_master_ruser),    //   input,    width = 8,                   .ruser
		.WUSER    (mgc_axi4_master_1_altera_axi4_master_wuser),    //  output,    width = 8,                   .wuser
		.RDATA    (mgc_axi4_master_1_altera_axi4_master_rdata),    //   input,  width = 256,                   .rdata
		.RID      (mgc_axi4_master_1_altera_axi4_master_rid),      //   input,    width = 7,                   .rid
		.WDATA    (mgc_axi4_master_1_altera_axi4_master_wdata),    //  output,  width = 256,                   .wdata
		.WSTRB    (mgc_axi4_master_1_altera_axi4_master_wstrb),    //  output,   width = 32,                   .wstrb
		.BID      (mgc_axi4_master_1_altera_axi4_master_bid),      //   input,    width = 7,                   .bid
		.ACLK     (iopll_0_outclk0_clk),                           //   input,    width = 1,         clock_sink.clk
		.ARESETn  (~rst_controller_reset_out_reset)                //   input,    width = 1,         reset_sink.reset_n
	);

	noc_reset noc_reset (
		.in_reset  (noc_reset_in_reset),        //   input,  width = 1,  in_reset.reset
		.out_reset (noc_reset_out_reset_reset)  //  output,  width = 1, out_reset.reset
	);

	my_sys_altera_mm_interconnect_1920_5ioayuq mm_interconnect_0 (
		.mgc_axi4_master_0_altera_axi4_master_awid                                             (mgc_axi4_master_0_altera_axi4_master_awid),               //   input,    width = 7,                                            mgc_axi4_master_0_altera_axi4_master.awid
		.mgc_axi4_master_0_altera_axi4_master_awaddr                                           (mgc_axi4_master_0_altera_axi4_master_awaddr),             //   input,   width = 64,                                                                                .awaddr
		.mgc_axi4_master_0_altera_axi4_master_awlen                                            (mgc_axi4_master_0_altera_axi4_master_awlen),              //   input,    width = 8,                                                                                .awlen
		.mgc_axi4_master_0_altera_axi4_master_awsize                                           (mgc_axi4_master_0_altera_axi4_master_awsize),             //   input,    width = 3,                                                                                .awsize
		.mgc_axi4_master_0_altera_axi4_master_awburst                                          (mgc_axi4_master_0_altera_axi4_master_awburst),            //   input,    width = 2,                                                                                .awburst
		.mgc_axi4_master_0_altera_axi4_master_awlock                                           (mgc_axi4_master_0_altera_axi4_master_awlock),             //   input,    width = 1,                                                                                .awlock
		.mgc_axi4_master_0_altera_axi4_master_awprot                                           (mgc_axi4_master_0_altera_axi4_master_awprot),             //   input,    width = 3,                                                                                .awprot
		.mgc_axi4_master_0_altera_axi4_master_awuser                                           (mgc_axi4_master_0_altera_axi4_master_awuser),             //   input,    width = 8,                                                                                .awuser
		.mgc_axi4_master_0_altera_axi4_master_awqos                                            (mgc_axi4_master_0_altera_axi4_master_awqos),              //   input,    width = 4,                                                                                .awqos
		.mgc_axi4_master_0_altera_axi4_master_awregion                                         (mgc_axi4_master_0_altera_axi4_master_awregion),           //   input,    width = 4,                                                                                .awregion
		.mgc_axi4_master_0_altera_axi4_master_awvalid                                          (mgc_axi4_master_0_altera_axi4_master_awvalid),            //   input,    width = 1,                                                                                .awvalid
		.mgc_axi4_master_0_altera_axi4_master_awready                                          (mgc_axi4_master_0_altera_axi4_master_awready),            //  output,    width = 1,                                                                                .awready
		.mgc_axi4_master_0_altera_axi4_master_wdata                                            (mgc_axi4_master_0_altera_axi4_master_wdata),              //   input,  width = 256,                                                                                .wdata
		.mgc_axi4_master_0_altera_axi4_master_wstrb                                            (mgc_axi4_master_0_altera_axi4_master_wstrb),              //   input,   width = 32,                                                                                .wstrb
		.mgc_axi4_master_0_altera_axi4_master_wlast                                            (mgc_axi4_master_0_altera_axi4_master_wlast),              //   input,    width = 1,                                                                                .wlast
		.mgc_axi4_master_0_altera_axi4_master_wvalid                                           (mgc_axi4_master_0_altera_axi4_master_wvalid),             //   input,    width = 1,                                                                                .wvalid
		.mgc_axi4_master_0_altera_axi4_master_wuser                                            (mgc_axi4_master_0_altera_axi4_master_wuser),              //   input,    width = 8,                                                                                .wuser
		.mgc_axi4_master_0_altera_axi4_master_wready                                           (mgc_axi4_master_0_altera_axi4_master_wready),             //  output,    width = 1,                                                                                .wready
		.mgc_axi4_master_0_altera_axi4_master_bid                                              (mgc_axi4_master_0_altera_axi4_master_bid),                //  output,    width = 7,                                                                                .bid
		.mgc_axi4_master_0_altera_axi4_master_bresp                                            (mgc_axi4_master_0_altera_axi4_master_bresp),              //  output,    width = 2,                                                                                .bresp
		.mgc_axi4_master_0_altera_axi4_master_bvalid                                           (mgc_axi4_master_0_altera_axi4_master_bvalid),             //  output,    width = 1,                                                                                .bvalid
		.mgc_axi4_master_0_altera_axi4_master_bready                                           (mgc_axi4_master_0_altera_axi4_master_bready),             //   input,    width = 1,                                                                                .bready
		.mgc_axi4_master_0_altera_axi4_master_arid                                             (mgc_axi4_master_0_altera_axi4_master_arid),               //   input,    width = 7,                                                                                .arid
		.mgc_axi4_master_0_altera_axi4_master_araddr                                           (mgc_axi4_master_0_altera_axi4_master_araddr),             //   input,   width = 64,                                                                                .araddr
		.mgc_axi4_master_0_altera_axi4_master_arlen                                            (mgc_axi4_master_0_altera_axi4_master_arlen),              //   input,    width = 8,                                                                                .arlen
		.mgc_axi4_master_0_altera_axi4_master_arsize                                           (mgc_axi4_master_0_altera_axi4_master_arsize),             //   input,    width = 3,                                                                                .arsize
		.mgc_axi4_master_0_altera_axi4_master_arburst                                          (mgc_axi4_master_0_altera_axi4_master_arburst),            //   input,    width = 2,                                                                                .arburst
		.mgc_axi4_master_0_altera_axi4_master_arlock                                           (mgc_axi4_master_0_altera_axi4_master_arlock),             //   input,    width = 1,                                                                                .arlock
		.mgc_axi4_master_0_altera_axi4_master_arprot                                           (mgc_axi4_master_0_altera_axi4_master_arprot),             //   input,    width = 3,                                                                                .arprot
		.mgc_axi4_master_0_altera_axi4_master_aruser                                           (mgc_axi4_master_0_altera_axi4_master_aruser),             //   input,    width = 8,                                                                                .aruser
		.mgc_axi4_master_0_altera_axi4_master_arqos                                            (mgc_axi4_master_0_altera_axi4_master_arqos),              //   input,    width = 4,                                                                                .arqos
		.mgc_axi4_master_0_altera_axi4_master_arregion                                         (mgc_axi4_master_0_altera_axi4_master_arregion),           //   input,    width = 4,                                                                                .arregion
		.mgc_axi4_master_0_altera_axi4_master_arvalid                                          (mgc_axi4_master_0_altera_axi4_master_arvalid),            //   input,    width = 1,                                                                                .arvalid
		.mgc_axi4_master_0_altera_axi4_master_arready                                          (mgc_axi4_master_0_altera_axi4_master_arready),            //  output,    width = 1,                                                                                .arready
		.mgc_axi4_master_0_altera_axi4_master_rid                                              (mgc_axi4_master_0_altera_axi4_master_rid),                //  output,    width = 7,                                                                                .rid
		.mgc_axi4_master_0_altera_axi4_master_rdata                                            (mgc_axi4_master_0_altera_axi4_master_rdata),              //  output,  width = 256,                                                                                .rdata
		.mgc_axi4_master_0_altera_axi4_master_rresp                                            (mgc_axi4_master_0_altera_axi4_master_rresp),              //  output,    width = 2,                                                                                .rresp
		.mgc_axi4_master_0_altera_axi4_master_rlast                                            (mgc_axi4_master_0_altera_axi4_master_rlast),              //  output,    width = 1,                                                                                .rlast
		.mgc_axi4_master_0_altera_axi4_master_rvalid                                           (mgc_axi4_master_0_altera_axi4_master_rvalid),             //  output,    width = 1,                                                                                .rvalid
		.mgc_axi4_master_0_altera_axi4_master_rready                                           (mgc_axi4_master_0_altera_axi4_master_rready),             //   input,    width = 1,                                                                                .rready
		.mgc_axi4_master_0_altera_axi4_master_ruser                                            (mgc_axi4_master_0_altera_axi4_master_ruser),              //  output,    width = 8,                                                                                .ruser
		.intel_noc_initiator_0_s0_axi4_awid                                                    (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awid),    //  output,    width = 7,                                                   intel_noc_initiator_0_s0_axi4.awid
		.intel_noc_initiator_0_s0_axi4_awaddr                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awaddr),  //  output,   width = 44,                                                                                .awaddr
		.intel_noc_initiator_0_s0_axi4_awlen                                                   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awlen),   //  output,    width = 8,                                                                                .awlen
		.intel_noc_initiator_0_s0_axi4_awsize                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awsize),  //  output,    width = 3,                                                                                .awsize
		.intel_noc_initiator_0_s0_axi4_awburst                                                 (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awburst), //  output,    width = 2,                                                                                .awburst
		.intel_noc_initiator_0_s0_axi4_awlock                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awlock),  //  output,    width = 1,                                                                                .awlock
		.intel_noc_initiator_0_s0_axi4_awprot                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awprot),  //  output,    width = 3,                                                                                .awprot
		.intel_noc_initiator_0_s0_axi4_awuser                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awuser),  //  output,   width = 11,                                                                                .awuser
		.intel_noc_initiator_0_s0_axi4_awqos                                                   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awqos),   //  output,    width = 4,                                                                                .awqos
		.intel_noc_initiator_0_s0_axi4_awvalid                                                 (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awvalid), //  output,    width = 1,                                                                                .awvalid
		.intel_noc_initiator_0_s0_axi4_awready                                                 (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_awready), //   input,    width = 1,                                                                                .awready
		.intel_noc_initiator_0_s0_axi4_wdata                                                   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wdata),   //  output,  width = 256,                                                                                .wdata
		.intel_noc_initiator_0_s0_axi4_wstrb                                                   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wstrb),   //  output,   width = 32,                                                                                .wstrb
		.intel_noc_initiator_0_s0_axi4_wlast                                                   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wlast),   //  output,    width = 1,                                                                                .wlast
		.intel_noc_initiator_0_s0_axi4_wvalid                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wvalid),  //  output,    width = 1,                                                                                .wvalid
		.intel_noc_initiator_0_s0_axi4_wuser                                                   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wuser),   //  output,   width = 32,                                                                                .wuser
		.intel_noc_initiator_0_s0_axi4_wready                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_wready),  //   input,    width = 1,                                                                                .wready
		.intel_noc_initiator_0_s0_axi4_bid                                                     (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_bid),     //   input,    width = 7,                                                                                .bid
		.intel_noc_initiator_0_s0_axi4_bresp                                                   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_bresp),   //   input,    width = 2,                                                                                .bresp
		.intel_noc_initiator_0_s0_axi4_bvalid                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_bvalid),  //   input,    width = 1,                                                                                .bvalid
		.intel_noc_initiator_0_s0_axi4_bready                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_bready),  //  output,    width = 1,                                                                                .bready
		.intel_noc_initiator_0_s0_axi4_arid                                                    (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arid),    //  output,    width = 7,                                                                                .arid
		.intel_noc_initiator_0_s0_axi4_araddr                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_araddr),  //  output,   width = 44,                                                                                .araddr
		.intel_noc_initiator_0_s0_axi4_arlen                                                   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arlen),   //  output,    width = 8,                                                                                .arlen
		.intel_noc_initiator_0_s0_axi4_arsize                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arsize),  //  output,    width = 3,                                                                                .arsize
		.intel_noc_initiator_0_s0_axi4_arburst                                                 (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arburst), //  output,    width = 2,                                                                                .arburst
		.intel_noc_initiator_0_s0_axi4_arlock                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arlock),  //  output,    width = 1,                                                                                .arlock
		.intel_noc_initiator_0_s0_axi4_arprot                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arprot),  //  output,    width = 3,                                                                                .arprot
		.intel_noc_initiator_0_s0_axi4_aruser                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_aruser),  //  output,   width = 11,                                                                                .aruser
		.intel_noc_initiator_0_s0_axi4_arqos                                                   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arqos),   //  output,    width = 4,                                                                                .arqos
		.intel_noc_initiator_0_s0_axi4_arvalid                                                 (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arvalid), //  output,    width = 1,                                                                                .arvalid
		.intel_noc_initiator_0_s0_axi4_arready                                                 (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_arready), //   input,    width = 1,                                                                                .arready
		.intel_noc_initiator_0_s0_axi4_rid                                                     (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rid),     //   input,    width = 7,                                                                                .rid
		.intel_noc_initiator_0_s0_axi4_rdata                                                   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rdata),   //   input,  width = 256,                                                                                .rdata
		.intel_noc_initiator_0_s0_axi4_rresp                                                   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rresp),   //   input,    width = 2,                                                                                .rresp
		.intel_noc_initiator_0_s0_axi4_rlast                                                   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rlast),   //   input,    width = 1,                                                                                .rlast
		.intel_noc_initiator_0_s0_axi4_rvalid                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rvalid),  //   input,    width = 1,                                                                                .rvalid
		.intel_noc_initiator_0_s0_axi4_rready                                                  (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_rready),  //  output,    width = 1,                                                                                .rready
		.intel_noc_initiator_0_s0_axi4_ruser                                                   (mm_interconnect_0_intel_noc_initiator_0_s0_axi4_ruser),   //   input,   width = 32,                                                                                .ruser
		.mgc_axi4_master_0_altera_axi4_master_translator_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                      //   input,    width = 1, mgc_axi4_master_0_altera_axi4_master_translator_clk_reset_reset_bridge_in_reset.reset
		.intel_noc_initiator_0_s0_axi4_translator_clk_reset_reset_bridge_in_reset_reset        (rst_controller_002_reset_out_reset),                      //   input,    width = 1,        intel_noc_initiator_0_s0_axi4_translator_clk_reset_reset_bridge_in_reset.reset
		.iopll_0_outclk0_clk                                                                   (iopll_0_outclk0_clk)                                      //   input,    width = 1,                                                                 iopll_0_outclk0.clk
	);

	my_sys_altera_mm_interconnect_1920_dxipmqi mm_interconnect_1 (
		.mgc_axi4_master_1_altera_axi4_master_awid                                             (mgc_axi4_master_1_altera_axi4_master_awid),               //   input,    width = 7,                                            mgc_axi4_master_1_altera_axi4_master.awid
		.mgc_axi4_master_1_altera_axi4_master_awaddr                                           (mgc_axi4_master_1_altera_axi4_master_awaddr),             //   input,   width = 64,                                                                                .awaddr
		.mgc_axi4_master_1_altera_axi4_master_awlen                                            (mgc_axi4_master_1_altera_axi4_master_awlen),              //   input,    width = 8,                                                                                .awlen
		.mgc_axi4_master_1_altera_axi4_master_awsize                                           (mgc_axi4_master_1_altera_axi4_master_awsize),             //   input,    width = 3,                                                                                .awsize
		.mgc_axi4_master_1_altera_axi4_master_awburst                                          (mgc_axi4_master_1_altera_axi4_master_awburst),            //   input,    width = 2,                                                                                .awburst
		.mgc_axi4_master_1_altera_axi4_master_awlock                                           (mgc_axi4_master_1_altera_axi4_master_awlock),             //   input,    width = 1,                                                                                .awlock
		.mgc_axi4_master_1_altera_axi4_master_awprot                                           (mgc_axi4_master_1_altera_axi4_master_awprot),             //   input,    width = 3,                                                                                .awprot
		.mgc_axi4_master_1_altera_axi4_master_awuser                                           (mgc_axi4_master_1_altera_axi4_master_awuser),             //   input,    width = 8,                                                                                .awuser
		.mgc_axi4_master_1_altera_axi4_master_awqos                                            (mgc_axi4_master_1_altera_axi4_master_awqos),              //   input,    width = 4,                                                                                .awqos
		.mgc_axi4_master_1_altera_axi4_master_awregion                                         (mgc_axi4_master_1_altera_axi4_master_awregion),           //   input,    width = 4,                                                                                .awregion
		.mgc_axi4_master_1_altera_axi4_master_awvalid                                          (mgc_axi4_master_1_altera_axi4_master_awvalid),            //   input,    width = 1,                                                                                .awvalid
		.mgc_axi4_master_1_altera_axi4_master_awready                                          (mgc_axi4_master_1_altera_axi4_master_awready),            //  output,    width = 1,                                                                                .awready
		.mgc_axi4_master_1_altera_axi4_master_wdata                                            (mgc_axi4_master_1_altera_axi4_master_wdata),              //   input,  width = 256,                                                                                .wdata
		.mgc_axi4_master_1_altera_axi4_master_wstrb                                            (mgc_axi4_master_1_altera_axi4_master_wstrb),              //   input,   width = 32,                                                                                .wstrb
		.mgc_axi4_master_1_altera_axi4_master_wlast                                            (mgc_axi4_master_1_altera_axi4_master_wlast),              //   input,    width = 1,                                                                                .wlast
		.mgc_axi4_master_1_altera_axi4_master_wvalid                                           (mgc_axi4_master_1_altera_axi4_master_wvalid),             //   input,    width = 1,                                                                                .wvalid
		.mgc_axi4_master_1_altera_axi4_master_wuser                                            (mgc_axi4_master_1_altera_axi4_master_wuser),              //   input,    width = 8,                                                                                .wuser
		.mgc_axi4_master_1_altera_axi4_master_wready                                           (mgc_axi4_master_1_altera_axi4_master_wready),             //  output,    width = 1,                                                                                .wready
		.mgc_axi4_master_1_altera_axi4_master_bid                                              (mgc_axi4_master_1_altera_axi4_master_bid),                //  output,    width = 7,                                                                                .bid
		.mgc_axi4_master_1_altera_axi4_master_bresp                                            (mgc_axi4_master_1_altera_axi4_master_bresp),              //  output,    width = 2,                                                                                .bresp
		.mgc_axi4_master_1_altera_axi4_master_bvalid                                           (mgc_axi4_master_1_altera_axi4_master_bvalid),             //  output,    width = 1,                                                                                .bvalid
		.mgc_axi4_master_1_altera_axi4_master_bready                                           (mgc_axi4_master_1_altera_axi4_master_bready),             //   input,    width = 1,                                                                                .bready
		.mgc_axi4_master_1_altera_axi4_master_arid                                             (mgc_axi4_master_1_altera_axi4_master_arid),               //   input,    width = 7,                                                                                .arid
		.mgc_axi4_master_1_altera_axi4_master_araddr                                           (mgc_axi4_master_1_altera_axi4_master_araddr),             //   input,   width = 64,                                                                                .araddr
		.mgc_axi4_master_1_altera_axi4_master_arlen                                            (mgc_axi4_master_1_altera_axi4_master_arlen),              //   input,    width = 8,                                                                                .arlen
		.mgc_axi4_master_1_altera_axi4_master_arsize                                           (mgc_axi4_master_1_altera_axi4_master_arsize),             //   input,    width = 3,                                                                                .arsize
		.mgc_axi4_master_1_altera_axi4_master_arburst                                          (mgc_axi4_master_1_altera_axi4_master_arburst),            //   input,    width = 2,                                                                                .arburst
		.mgc_axi4_master_1_altera_axi4_master_arlock                                           (mgc_axi4_master_1_altera_axi4_master_arlock),             //   input,    width = 1,                                                                                .arlock
		.mgc_axi4_master_1_altera_axi4_master_arprot                                           (mgc_axi4_master_1_altera_axi4_master_arprot),             //   input,    width = 3,                                                                                .arprot
		.mgc_axi4_master_1_altera_axi4_master_aruser                                           (mgc_axi4_master_1_altera_axi4_master_aruser),             //   input,    width = 8,                                                                                .aruser
		.mgc_axi4_master_1_altera_axi4_master_arqos                                            (mgc_axi4_master_1_altera_axi4_master_arqos),              //   input,    width = 4,                                                                                .arqos
		.mgc_axi4_master_1_altera_axi4_master_arregion                                         (mgc_axi4_master_1_altera_axi4_master_arregion),           //   input,    width = 4,                                                                                .arregion
		.mgc_axi4_master_1_altera_axi4_master_arvalid                                          (mgc_axi4_master_1_altera_axi4_master_arvalid),            //   input,    width = 1,                                                                                .arvalid
		.mgc_axi4_master_1_altera_axi4_master_arready                                          (mgc_axi4_master_1_altera_axi4_master_arready),            //  output,    width = 1,                                                                                .arready
		.mgc_axi4_master_1_altera_axi4_master_rid                                              (mgc_axi4_master_1_altera_axi4_master_rid),                //  output,    width = 7,                                                                                .rid
		.mgc_axi4_master_1_altera_axi4_master_rdata                                            (mgc_axi4_master_1_altera_axi4_master_rdata),              //  output,  width = 256,                                                                                .rdata
		.mgc_axi4_master_1_altera_axi4_master_rresp                                            (mgc_axi4_master_1_altera_axi4_master_rresp),              //  output,    width = 2,                                                                                .rresp
		.mgc_axi4_master_1_altera_axi4_master_rlast                                            (mgc_axi4_master_1_altera_axi4_master_rlast),              //  output,    width = 1,                                                                                .rlast
		.mgc_axi4_master_1_altera_axi4_master_rvalid                                           (mgc_axi4_master_1_altera_axi4_master_rvalid),             //  output,    width = 1,                                                                                .rvalid
		.mgc_axi4_master_1_altera_axi4_master_rready                                           (mgc_axi4_master_1_altera_axi4_master_rready),             //   input,    width = 1,                                                                                .rready
		.mgc_axi4_master_1_altera_axi4_master_ruser                                            (mgc_axi4_master_1_altera_axi4_master_ruser),              //  output,    width = 8,                                                                                .ruser
		.intel_noc_initiator_0_s1_axi4_awid                                                    (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awid),    //  output,    width = 7,                                                   intel_noc_initiator_0_s1_axi4.awid
		.intel_noc_initiator_0_s1_axi4_awaddr                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awaddr),  //  output,   width = 44,                                                                                .awaddr
		.intel_noc_initiator_0_s1_axi4_awlen                                                   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awlen),   //  output,    width = 8,                                                                                .awlen
		.intel_noc_initiator_0_s1_axi4_awsize                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awsize),  //  output,    width = 3,                                                                                .awsize
		.intel_noc_initiator_0_s1_axi4_awburst                                                 (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awburst), //  output,    width = 2,                                                                                .awburst
		.intel_noc_initiator_0_s1_axi4_awlock                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awlock),  //  output,    width = 1,                                                                                .awlock
		.intel_noc_initiator_0_s1_axi4_awprot                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awprot),  //  output,    width = 3,                                                                                .awprot
		.intel_noc_initiator_0_s1_axi4_awuser                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awuser),  //  output,   width = 11,                                                                                .awuser
		.intel_noc_initiator_0_s1_axi4_awqos                                                   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awqos),   //  output,    width = 4,                                                                                .awqos
		.intel_noc_initiator_0_s1_axi4_awvalid                                                 (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awvalid), //  output,    width = 1,                                                                                .awvalid
		.intel_noc_initiator_0_s1_axi4_awready                                                 (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_awready), //   input,    width = 1,                                                                                .awready
		.intel_noc_initiator_0_s1_axi4_wdata                                                   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wdata),   //  output,  width = 256,                                                                                .wdata
		.intel_noc_initiator_0_s1_axi4_wstrb                                                   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wstrb),   //  output,   width = 32,                                                                                .wstrb
		.intel_noc_initiator_0_s1_axi4_wlast                                                   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wlast),   //  output,    width = 1,                                                                                .wlast
		.intel_noc_initiator_0_s1_axi4_wvalid                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wvalid),  //  output,    width = 1,                                                                                .wvalid
		.intel_noc_initiator_0_s1_axi4_wuser                                                   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wuser),   //  output,   width = 32,                                                                                .wuser
		.intel_noc_initiator_0_s1_axi4_wready                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_wready),  //   input,    width = 1,                                                                                .wready
		.intel_noc_initiator_0_s1_axi4_bid                                                     (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_bid),     //   input,    width = 7,                                                                                .bid
		.intel_noc_initiator_0_s1_axi4_bresp                                                   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_bresp),   //   input,    width = 2,                                                                                .bresp
		.intel_noc_initiator_0_s1_axi4_bvalid                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_bvalid),  //   input,    width = 1,                                                                                .bvalid
		.intel_noc_initiator_0_s1_axi4_bready                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_bready),  //  output,    width = 1,                                                                                .bready
		.intel_noc_initiator_0_s1_axi4_arid                                                    (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arid),    //  output,    width = 7,                                                                                .arid
		.intel_noc_initiator_0_s1_axi4_araddr                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_araddr),  //  output,   width = 44,                                                                                .araddr
		.intel_noc_initiator_0_s1_axi4_arlen                                                   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arlen),   //  output,    width = 8,                                                                                .arlen
		.intel_noc_initiator_0_s1_axi4_arsize                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arsize),  //  output,    width = 3,                                                                                .arsize
		.intel_noc_initiator_0_s1_axi4_arburst                                                 (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arburst), //  output,    width = 2,                                                                                .arburst
		.intel_noc_initiator_0_s1_axi4_arlock                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arlock),  //  output,    width = 1,                                                                                .arlock
		.intel_noc_initiator_0_s1_axi4_arprot                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arprot),  //  output,    width = 3,                                                                                .arprot
		.intel_noc_initiator_0_s1_axi4_aruser                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_aruser),  //  output,   width = 11,                                                                                .aruser
		.intel_noc_initiator_0_s1_axi4_arqos                                                   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arqos),   //  output,    width = 4,                                                                                .arqos
		.intel_noc_initiator_0_s1_axi4_arvalid                                                 (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arvalid), //  output,    width = 1,                                                                                .arvalid
		.intel_noc_initiator_0_s1_axi4_arready                                                 (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_arready), //   input,    width = 1,                                                                                .arready
		.intel_noc_initiator_0_s1_axi4_rid                                                     (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rid),     //   input,    width = 7,                                                                                .rid
		.intel_noc_initiator_0_s1_axi4_rdata                                                   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rdata),   //   input,  width = 256,                                                                                .rdata
		.intel_noc_initiator_0_s1_axi4_rresp                                                   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rresp),   //   input,    width = 2,                                                                                .rresp
		.intel_noc_initiator_0_s1_axi4_rlast                                                   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rlast),   //   input,    width = 1,                                                                                .rlast
		.intel_noc_initiator_0_s1_axi4_rvalid                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rvalid),  //   input,    width = 1,                                                                                .rvalid
		.intel_noc_initiator_0_s1_axi4_rready                                                  (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_rready),  //  output,    width = 1,                                                                                .rready
		.intel_noc_initiator_0_s1_axi4_ruser                                                   (mm_interconnect_1_intel_noc_initiator_0_s1_axi4_ruser),   //   input,   width = 32,                                                                                .ruser
		.mgc_axi4_master_1_altera_axi4_master_translator_clk_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                      //   input,    width = 1, mgc_axi4_master_1_altera_axi4_master_translator_clk_reset_reset_bridge_in_reset.reset
		.intel_noc_initiator_0_s1_axi4_translator_clk_reset_reset_bridge_in_reset_reset        (rst_controller_002_reset_out_reset),                      //   input,    width = 1,        intel_noc_initiator_0_s1_axi4_translator_clk_reset_reset_bridge_in_reset.reset
		.iopll_0_outclk0_clk                                                                   (iopll_0_outclk0_clk)                                      //   input,    width = 1,                                                                 iopll_0_outclk0.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (axi_reset_out_reset_reset),      //   input,  width = 1, reset_in0.reset
		.clk            (iopll_0_outclk0_clk),            //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                               // (terminated),                       
		.reset_req_in0  (1'b0),                           // (terminated),                       
		.reset_in1      (1'b0),                           // (terminated),                       
		.reset_req_in1  (1'b0),                           // (terminated),                       
		.reset_in2      (1'b0),                           // (terminated),                       
		.reset_req_in2  (1'b0),                           // (terminated),                       
		.reset_in3      (1'b0),                           // (terminated),                       
		.reset_req_in3  (1'b0),                           // (terminated),                       
		.reset_in4      (1'b0),                           // (terminated),                       
		.reset_req_in4  (1'b0),                           // (terminated),                       
		.reset_in5      (1'b0),                           // (terminated),                       
		.reset_req_in5  (1'b0),                           // (terminated),                       
		.reset_in6      (1'b0),                           // (terminated),                       
		.reset_req_in6  (1'b0),                           // (terminated),                       
		.reset_in7      (1'b0),                           // (terminated),                       
		.reset_req_in7  (1'b0),                           // (terminated),                       
		.reset_in8      (1'b0),                           // (terminated),                       
		.reset_req_in8  (1'b0),                           // (terminated),                       
		.reset_in9      (1'b0),                           // (terminated),                       
		.reset_req_in9  (1'b0),                           // (terminated),                       
		.reset_in10     (1'b0),                           // (terminated),                       
		.reset_req_in10 (1'b0),                           // (terminated),                       
		.reset_in11     (1'b0),                           // (terminated),                       
		.reset_req_in11 (1'b0),                           // (terminated),                       
		.reset_in12     (1'b0),                           // (terminated),                       
		.reset_req_in12 (1'b0),                           // (terminated),                       
		.reset_in13     (1'b0),                           // (terminated),                       
		.reset_req_in13 (1'b0),                           // (terminated),                       
		.reset_in14     (1'b0),                           // (terminated),                       
		.reset_req_in14 (1'b0),                           // (terminated),                       
		.reset_in15     (1'b0),                           // (terminated),                       
		.reset_req_in15 (1'b0)                            // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (axi_reset_out_reset_reset),          //   input,  width = 1, reset_in0.reset
		.clk            (iopll_0_outclk0_clk),                //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (noc_reset_out_reset_reset),          //   input,  width = 1, reset_in0.reset
		.clk            (iopll_0_outclk0_clk),                //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule
